/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 */
class add_test extends random_test;
    `uvm_component_utils(add_test)

//------------------------------------------------------------------------------
// local variables
//------------------------------------------------------------------------------
  //  env env_h;

//------------------------------------------------------------------------------
// constructor
//------------------------------------------------------------------------------
    function new (string name, uvm_component parent);
        super.new(name,parent);
    endfunction : new

//------------------------------------------------------------------------------
// build phase
//------------------------------------------------------------------------------

      function void build_phase(uvm_phase phase);
        
        super.build_phase(phase);

        // set the factory to produce a corner_tpgen whenever it would produce
        // a random_tpgen
        random_tpgen::type_id::set_type_override(corners_tpgen::get_type());

    endfunction : build_phase

endclass


